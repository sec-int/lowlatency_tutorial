//////////////////////////////////////////////////
// mixt module
//
module  mixt  ( a , y ) ;


input    [0:63]  a  ;

output   [0:63]  y  ;

wire     [0:63]  coef1  [0:63] ;

// Matrix definitions
//
assign  coef1[00] = 64'b0000100010001000000000000000000000000000000000000000000000000000 ;
assign  coef1[01] = 64'b0100000001000100000000000000000000000000000000000000000000000000 ;
assign  coef1[02] = 64'b0010001000000010000000000000000000000000000000000000000000000000 ;
assign  coef1[03] = 64'b0001000100010000000000000000000000000000000000000000000000000000 ;
assign  coef1[04] = 64'b1000100010000000000000000000000000000000000000000000000000000000 ;
assign  coef1[05] = 64'b0000010001000100000000000000000000000000000000000000000000000000 ;
assign  coef1[06] = 64'b0010000000100010000000000000000000000000000000000000000000000000 ;
assign  coef1[07] = 64'b0001000100000001000000000000000000000000000000000000000000000000 ;
assign  coef1[08] = 64'b1000100000001000000000000000000000000000000000000000000000000000 ;
assign  coef1[09] = 64'b0100010001000000000000000000000000000000000000000000000000000000 ;
assign  coef1[10] = 64'b0000001000100010000000000000000000000000000000000000000000000000 ;
assign  coef1[11] = 64'b0001000000010001000000000000000000000000000000000000000000000000 ;
assign  coef1[12] = 64'b1000000010001000000000000000000000000000000000000000000000000000 ;
assign  coef1[13] = 64'b0100010000000100000000000000000000000000000000000000000000000000 ;
assign  coef1[14] = 64'b0010001000100000000000000000000000000000000000000000000000000000 ;
assign  coef1[15] = 64'b0000000100010001000000000000000000000000000000000000000000000000 ;
assign  coef1[16] = 64'b0000000000000000100010001000000000000000000000000000000000000000 ;
assign  coef1[17] = 64'b0000000000000000000001000100010000000000000000000000000000000000 ;
assign  coef1[18] = 64'b0000000000000000001000000010001000000000000000000000000000000000 ;
assign  coef1[19] = 64'b0000000000000000000100010000000100000000000000000000000000000000 ;
assign  coef1[20] = 64'b0000000000000000100010000000100000000000000000000000000000000000 ;
assign  coef1[21] = 64'b0000000000000000010001000100000000000000000000000000000000000000 ;
assign  coef1[22] = 64'b0000000000000000000000100010001000000000000000000000000000000000 ;
assign  coef1[23] = 64'b0000000000000000000100000001000100000000000000000000000000000000 ;
assign  coef1[24] = 64'b0000000000000000100000001000100000000000000000000000000000000000 ;
assign  coef1[25] = 64'b0000000000000000010001000000010000000000000000000000000000000000 ;
assign  coef1[26] = 64'b0000000000000000001000100010000000000000000000000000000000000000 ;
assign  coef1[27] = 64'b0000000000000000000000010001000100000000000000000000000000000000 ;
assign  coef1[28] = 64'b0000000000000000000010001000100000000000000000000000000000000000 ;
assign  coef1[29] = 64'b0000000000000000010000000100010000000000000000000000000000000000 ;
assign  coef1[30] = 64'b0000000000000000001000100000001000000000000000000000000000000000 ;
assign  coef1[31] = 64'b0000000000000000000100010001000000000000000000000000000000000000 ;
assign  coef1[32] = 64'b0000000000000000000000000000000010001000100000000000000000000000 ;
assign  coef1[33] = 64'b0000000000000000000000000000000000000100010001000000000000000000 ;
assign  coef1[34] = 64'b0000000000000000000000000000000000100000001000100000000000000000 ;
assign  coef1[35] = 64'b0000000000000000000000000000000000010001000000010000000000000000 ;
assign  coef1[36] = 64'b0000000000000000000000000000000010001000000010000000000000000000 ;
assign  coef1[37] = 64'b0000000000000000000000000000000001000100010000000000000000000000 ;
assign  coef1[38] = 64'b0000000000000000000000000000000000000010001000100000000000000000 ;
assign  coef1[39] = 64'b0000000000000000000000000000000000010000000100010000000000000000 ;
assign  coef1[40] = 64'b0000000000000000000000000000000010000000100010000000000000000000 ;
assign  coef1[41] = 64'b0000000000000000000000000000000001000100000001000000000000000000 ;
assign  coef1[42] = 64'b0000000000000000000000000000000000100010001000000000000000000000 ;
assign  coef1[43] = 64'b0000000000000000000000000000000000000001000100010000000000000000 ;
assign  coef1[44] = 64'b0000000000000000000000000000000000001000100010000000000000000000 ;
assign  coef1[45] = 64'b0000000000000000000000000000000001000000010001000000000000000000 ;
assign  coef1[46] = 64'b0000000000000000000000000000000000100010000000100000000000000000 ;
assign  coef1[47] = 64'b0000000000000000000000000000000000010001000100000000000000000000 ;
assign  coef1[48] = 64'b0000000000000000000000000000000000000000000000000000100010001000 ;
assign  coef1[49] = 64'b0000000000000000000000000000000000000000000000000100000001000100 ;
assign  coef1[50] = 64'b0000000000000000000000000000000000000000000000000010001000000010 ;
assign  coef1[51] = 64'b0000000000000000000000000000000000000000000000000001000100010000 ;
assign  coef1[52] = 64'b0000000000000000000000000000000000000000000000001000100010000000 ;
assign  coef1[53] = 64'b0000000000000000000000000000000000000000000000000000010001000100 ;
assign  coef1[54] = 64'b0000000000000000000000000000000000000000000000000010000000100010 ;
assign  coef1[55] = 64'b0000000000000000000000000000000000000000000000000001000100000001 ;
assign  coef1[56] = 64'b0000000000000000000000000000000000000000000000001000100000001000 ;
assign  coef1[57] = 64'b0000000000000000000000000000000000000000000000000100010001000000 ;
assign  coef1[58] = 64'b0000000000000000000000000000000000000000000000000000001000100010 ;
assign  coef1[59] = 64'b0000000000000000000000000000000000000000000000000001000000010001 ;
assign  coef1[60] = 64'b0000000000000000000000000000000000000000000000001000000010001000 ;
assign  coef1[61] = 64'b0000000000000000000000000000000000000000000000000100010000000100 ;
assign  coef1[62] = 64'b0000000000000000000000000000000000000000000000000010001000100000 ;
assign  coef1[63] = 64'b0000000000000000000000000000000000000000000000000000000100010001 ;

// Multiply
//
genvar  i ;
generate
  for  ( i  =  0 ;  i  <  64 ;  i  =  i + 1 )
    begin  :  mixt
       assign  y[i] = ^ ( a & coef1[i] ) ;      
    end
endgenerate


endmodule

